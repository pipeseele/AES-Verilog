`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.01.2024 16:36:15
// Design Name: 
// Module Name: mul_2_module
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module gf256mult(a, b, z);
input [7:0] a;
input [7:0] b;
output [7:0] z;

assign z[0] = b[0]&a[0]^b[1]&a[7]^b[7]&a[1]^b[2]&a[6]^b[6]&a[2]^b[3]&a[5]^b[5]&a[3]^b[4]&a[4]^b[5]&a[7]^b[7]&a[5]^b[6]&a[6]^b[6]&a[7]^b[7]&a[6];

assign z[1] = b[0]&a[1]^b[1]&a[0]^b[1]&a[7]^b[7]&a[1]^b[2]&a[6]^b[6]&a[2]^b[2]&a[7]^b[7]&a[2]^b[3]&a[5]^b[5]&a[3]^b[3]&a[6]^b[6]&a[3]^b[4]&a[4]^b[4]&a[5]^b[5]&a[4]^b[5]&a[7]^b[7]&a[5]^b[6]&a[6]^b[7]&a[7];

assign z[2] = b[0]&a[2]^b[2]&a[0]^b[1]&a[1]^b[2]&a[7]^b[7]&a[2]^b[3]&a[6]^b[6]&a[3]^b[3]&a[7]^b[7]&a[3]^b[4]&a[5]^b[5]&a[4]^b[4]&a[6]^b[6]&a[4]^b[5]&a[5]^b[6]&a[7]^b[7]&a[6];

assign z[3] = b[0]&a[3]^b[3]&a[0]^b[1]&a[2]^b[2]&a[1]^b[1]&a[7]^b[7]&a[1]^b[2]&a[6]^b[6]&a[2]^b[3]&a[5]^b[5]&a[3]^b[3]&a[7]^b[7]&a[3]^b[4]&a[4]^b[4]&a[6]^b[6]&a[4]^b[4]&a[7]^b[7]&a[4]^b[5]&a[5]^b[5]&a[6]^b[6]&a[5]^b[5]&a[7]^b[7]&a[5]^b[6]&a[6]^b[6]&a[7]^b[7]&a[6]^b[7]&a[7];

assign z[4] = b[0]&a[4]^b[4]&a[0]^b[1]&a[3]^b[3]&a[1]^b[1]&a[7]^b[7]&a[1]^b[2]&a[2]^b[2]&a[6]^b[6]&a[2]^b[2]&a[7]^b[7]&a[2]^b[3]&a[5]^b[5]&a[3]^b[3]&a[6]^b[6]&a[3]^b[4]&a[4]^b[4]&a[5]^b[5]&a[4]^b[4]&a[7]^b[7]&a[4]^b[5]&a[6]^b[6]&a[5]^b[7]&a[7];

assign z[5] = b[0]&a[5]^b[5]&a[0]^b[1]&a[4]^b[4]&a[1]^b[2]&a[3]^b[3]&a[2]^b[2]&a[7]^b[7]&a[2]^b[3]&a[6]^b[6]&a[3]^b[3]&a[7]^b[7]&a[3]^b[4]&a[5]^b[5]&a[4]^b[4]&a[6]^b[6]&a[4]^b[5]&a[5]^b[5]&a[7]^b[7]&a[5]^b[6]&a[6];

assign z[6] = b[0]&a[6]^b[6]&a[0]^b[1]&a[5]^b[5]&a[1]^b[2]&a[4]^b[4]&a[2]^b[3]&a[3]^b[3]&a[7]^b[7]&a[3]^b[4]&a[6]^b[6]&a[4]^b[4]&a[7]^b[7]&a[4]^b[5]&a[5]^b[5]&a[6]^b[6]&a[5]^b[6]&a[7]^b[7]&a[6];

assign z[7] = b[0]&a[7]^b[7]&a[0]^b[1]&a[6]^b[6]&a[1]^b[2]&a[5]^b[5]&a[2]^b[3]&a[4]^b[4]&a[3]^b[4]&a[7]^b[7]&a[4]^b[5]&a[6]^b[6]&a[5]^b[5]&a[7]^b[7]&a[5]^b[6]&a[6]^b[7]&a[7];

endmodule